library ieee;
use ieee.std_logic_1164.all;
use work.common.all;

entity cpu is

end cpu;

architecture arch of cpu is
begin

end arch;

